library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity main is
end main;

architecture Behavioral of main is

begin


end Behavioral;

